`timescale 1ns / 1ps
//-------------------------------------------------------------------------------------------


//端口定义------------------------------------------------------------------------------------
module D_Splitter(
    input [31:0] Instr,
    output [5:0] D_opcode,
    output [4:0] D_rs,
    output [4:0] D_rt,
    output [4:0] D_rd,
    output [5:0] D_func,
    output [15:0] D_imm16,
    output [25:0] D_imm26
    );
//---------------------------------------------------------------------------------------------


//splitter-------------------------------------------------------------------------------------
    assign D_opcode = Instr[31:26];
    assign D_rs = Instr[25:21];
    assign D_rt = Instr[20:16];
    assign D_rd = Instr[15:11];
    assign D_func = Instr[5:0];
    assign D_imm16 = Instr[15:0];
    assign D_imm26 = Instr[25:0];
//----------------------------------------------------------------------------------------------

endmodule