`timescale 1ns / 1ps
//-----------------------------------------------------------------------------------------------------------------


//端口定义--------------------------------------------------------------------------------------------------------
module D_CMP (
    input [31:0] rs_Data,
    input [31:0] rt_Data,
    input [1:0] CU_CMP_op,
    output D_CMP_out
    );
//--------------------------------------------------------------------------------------------------------------    


//----------------------------------------------------------------------------------------------------------------
    assign D_CMP_out = (CU_CMP_op == 2'b01) ? (rs_Data != rt_Data) : 
                                             (rs_Data == rt_Data);
//---------------------------------------------------------------------------------------------------------------

endmodule