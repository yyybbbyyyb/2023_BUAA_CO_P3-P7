`timescale 1ns / 1ps
//-----------------------------------------------------------------------------
`define aluAdd    4'b0000
`define aluSub    4'b0001
`define aluOr     4'b0010
`define aluAnd    4'b0011
`define aluLui    4'b0100
//-------------------------------------------------------------------------------


//端口定义------------------------------------------------------------------------
module E_ALU(
    input [31:0] ALU_a,
    input [31:0] ALU_b,
    input [3:0] CU_ALU_op,
    output [31:0] E_ALU_out
    );
//---------------------------------------------------------------------------------	
      

//select_area----------------------------------------------------------------------    
    assign E_ALU_out = (CU_ALU_op == `aluAdd) ? ALU_a + ALU_b :           //加运�
                     (CU_ALU_op == `aluSub) ? ALU_a - ALU_b :           //减运�
                     (CU_ALU_op == `aluOr) ? ALU_a | ALU_b :            //或运�
                     (CU_ALU_op == `aluAnd) ? ALU_a & ALU_b :           //和运�
                     (CU_ALU_op == `aluLui) ? {ALU_b[15:0], 16'H0000} : //�6位补0
                     32'H0000_0000;
//----------------------------------------------------------------------------------


endmodule
