`timescale 1ns / 1ps
//-------------------------------------------------------------------------------------------


//端口定义--------------------------------------------------------------------------------------------------------
module F_D (
    input clk,
    input reset,
    input HCU_EN_FD,
    input HCU_clr_FD,
    input [31:0] F_Instr,
    input [31:0] F_PC,
    output reg [31:0] D_Instr,
    output reg [31:0] D_PC
    );
//----------------------------------------------------------------------------------------------------


//D_reg-------------------------------------------------------------------------------------------
    always @(posedge clk) begin
        if (reset | HCU_clr_FD) begin
            D_Instr <= 32'H0000_0000;
            D_PC <= 32'H0000_0000;
        end
        else begin
            if (HCU_EN_FD) begin
                D_Instr <= F_Instr;
                D_PC <= F_PC;
            end
        end
    end
//--------------------------------------------------------------------------------------------------


endmodule