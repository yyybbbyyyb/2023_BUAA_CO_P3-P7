`timescale 1ns / 1ps
//---------------------------------------------------------------------------------------------------------------------
`define dmWord    2'b00
`define dmByte    2'b01
`define dmHalf    2'b10
//--------------------------------------------------------------------------------------------------------------------


//端口定义--------------------------------------------------------------------------------------------------------------
module M_DMOUT (
    input [31:0] addr,            
    input [31:0] readData,
    input [1:0] CU_DM_op,
    input is_load,
    input is_addrOv,
    output reg [31:0] M_DM_out,
    output M_is_AdEL
    );
//---------------------------------------------------------------------------------------------------------------------------------
 
 
//define wire---------------------------------------------------------------------------------------------------------------------------
    wire [1:0] opB = addr[1:0];                             
    wire opHw = addr[1];                                     
    
    wire [7:0] B1 = readData[7:0];                   
    wire [7:0] B2 = readData[15:8];
    wire [7:0] B3 = readData[23:16];
    wire [7:0] B4 = readData[31:24];
    wire [15:0] Hw1 = readData[15:0];                 
    wire [15:0] Hw2 = readData[31:16];
//------------------------------------------------------------------------------------------------------------------------------------
  
  
//read-----------------------------------------------------------------------------------------------------------------------------------                                    
    always @(*) begin
        if (CU_DM_op == `dmWord) begin
            M_DM_out = readData;           
        end
        else if (CU_DM_op == `dmByte) begin
            case (opB)
                2'b00:  M_DM_out = {{24{B1[7]}}, B1};
                2'b01:  M_DM_out = {{24{B2[7]}}, B2};
                2'b10:  M_DM_out = {{24{B3[7]}}, B3};
                2'b11:  M_DM_out = {{24{B4[7]}}, B4};
            endcase
        end
        else if (CU_DM_op == `dmHalf) begin
            case (opHw)
                0:  M_DM_out = {{16{Hw1[15]}}, Hw1};
                1:  M_DM_out = {{16{Hw2[15]}}, Hw2};
            endcase
        end 
    end            
//-------------------------------------------------------------------------------------------------------------------------------


//exc_hand-------------------------------------------------------------------------------------------------------------------------------
    wire error_align = ((CU_DM_op == `dmWord) && (|addr[1:0])) ||
                       ((CU_DM_op == `dmHalf) && (addr[0]));
    
    wire error_outOfRange = !(((addr >= 32'H0000_0000) && (addr <= 32'H0000_2FFF)) ||
                              ((addr >= 32'H0000_7F00) && (addr <= 32'H0000_7F0B)) ||
                              ((addr >= 32'H0000_7F10) && (addr <= 32'H0000_7F1B)) ||
                              ((addr >= 32'H0000_7F20) && (addr <= 32'H0000_7F23)));
    
    wire error_timer = (CU_DM_op != `dmWord && 
                        (((addr >= 32'H0000_7F00) && (addr <= 32'H0000_7F0B)) ||
                         ((addr >= 32'H0000_7F10) && (addr <= 32'H0000_7F1B))));

    assign M_is_AdEL = (is_load) & (error_align | error_outOfRange | error_timer | is_addrOv);
//---------------------------------------------------------------------------------------------------------------------------------------
endmodule