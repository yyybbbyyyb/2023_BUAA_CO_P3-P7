`timescale 1ns / 1ps
//-----------------------------------------------------------------------------


//端口定义------------------------------------------------------------------------
module D_EXT (
    input [15:0] imm16,
    input CU_EXT_op,
    output [31:0] D_imm32
    );
//---------------------------------------------------------------------------------


//---------------------------------------------------------------------------------
    assign D_imm32 = (CU_EXT_op == 1) ? {{16{imm16[15]}}, imm16} :
                                        {16'H0000, imm16}; 
//----------------------------------------------------------------------------------


endmodule