`timescale 1ns / 1ps
//-----------------------------------------------------------------------------------------------------------------
`define npcPC4    3'b000
`define npcJal    3'b001
`define npcJr     3'b010
`define npcBranch 3'b011
`define npcEret   3'b100
//--------------------------------------------------------------------------------------------------------------


//端口定义-----------------------------------------------------------------------------------------------------
module D_NPC (
    input [31:0] F_PC,
    input [31:0] D_PC,   
    input [25:0] imm26,
    input [31:0] ra_Data,
    input CMP_out,
    input [2:0] CU_NPC_op,
    input req,
    input [31:0] EPC,
    output [31:0] NPC
    );
//------------------------------------------------------------------------------------------------


//select_area------------------------------------------------------------------------------------                 
    assign NPC = (req) ? 32'H0000_4180 :
                 (CU_NPC_op == `npcEret) ? EPC + 4 :   
                 (CU_NPC_op == `npcPC4) ? F_PC + 4 : 
                 (CU_NPC_op == `npcJal) ? {D_PC[31:28], imm26, 2'b00} :
                 (CU_NPC_op == `npcJr)  ? ra_Data :
                 (CU_NPC_op == `npcBranch && CMP_out) ? D_PC + 4 + {{14{imm26[15]}}, imm26[15:0], 2'b00} :
                 F_PC + 4;
//------------------------------------------------------------------------------------------------

endmodule