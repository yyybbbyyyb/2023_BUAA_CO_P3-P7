`timescale 1ns / 1ps
//-----------------------------------------------------------------------------------


//端口定义----------------------------------------------------------------------------
module F_IFU(
    input clk,
    input reset,
    input req,
    input HCU_EN_IFU,
    input [31:0] NPC,
    output reg [31:0] F_PC
    );
//-------------------------------------------------------------------------------------    


//初始化PC-----------------------------------------------------------------------------
    initial begin
        F_PC = 32'H0000_3000;
    end
//---------------------------------------------------------------------------------------


//PC-------------------------------------------------------------------------------------
    always @(posedge clk) begin
        if (reset) begin
            F_PC <= 32'H0000_3000;
        end
        else begin
            if (req) begin
                F_PC <= 32'H0000_4180;
            end
            else if (HCU_EN_IFU) begin
                F_PC <= NPC;        
            end
        end
    end
//-----------------------------------------------------------------------------------------

endmodule